// Copyright (c) 2012-2013 Ludvig Strigeus
// This program is GPL Licensed. See COPYING for the full license.

module TftDriver(input clk,
                 output reg tft_h, output reg tft_v,
                 output reg [3:0] tft_r, output reg[3:0] tft_g, output reg[3:0] tft_b,
                 input [14:0] pixel,        // Pixel for current cycle.
                 input de,
                 input border, output tft_clk);


endmodule

